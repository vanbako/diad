`ifndef SR_VH
`define SR_VH

`define INDEX_PC 0
`define INDEX_LR 1

`endif