`ifndef SR_VH
`define SR_VH

`define INDEX_FL  0
`define INDEX_LR  1
`define INDEX_IR  2
`define INDEX_SSP 3
`define INDEX_PC  0xf

`endif