`ifndef CC_VH
`define CC_VH

`define CC_RA 4'h0
`define CC_EQ 4'h1
`define CC_NE 4'h2
`define CC_LT 4'h3
`define CC_GT 4'h4
`define CC_LE 4'h5
`define CC_GE 4'h6

`endif
