`ifndef SIZES_VH
`define SIZES_VH

`define SIZE_ADDR 24
`define SIZE_DATA 24

`define HBIT_ADDR 23
`define HBIT_DATA 23

`endif
